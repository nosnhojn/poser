module module4 #(a bunch of stuff)(bar, foo);
  input bar;
  output foo;
endmodule
