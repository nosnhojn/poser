`include "this and"
`define this
module module0(bar, foo);
  input bar;
  output foo;
endmodule
