module module5(clk_, rst_, bar, foo);
  input clk_, rst_;
  input [1:0] bar;
  output foo;
endmodule
