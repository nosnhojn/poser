module poserCell
(
  clk,
  rst,
  i,
  o
);

parameter cellType = 0;
parameter activeRst = 0;

input clk;
input rst;
input i;
output o;

endmodule

