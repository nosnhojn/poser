module module5 (bar, foo);
  input bar;
  parameter blah ,a==,blah blah = llsdkfj,,;
  output foo;
endmodule
