module module1 (
  input bar,
  output foo
);
endmodule
