module module6(clk_, rst_, bar, foo);
  input clk_, rst_;
  input [1:0] bar;
  output [1:0] foo;
endmodule
