module module5(bar, foo);
  parameter blah ,a==,blah blah = llsdkfj,,;
  input bar;
  output foo;
endmodule
