module module0(clk, rst_n, bar, foo);
  input clk, rst_n;
  input [1:0] bar;
  output [1:0] foo;
endmodule
