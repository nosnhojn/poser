module module1(clk_, rst_, bar0, bar1, foo0, foo1);
  input clk_, rst_;
  input [1:0] bar0;
  input [1:0] bar1;
  output [1:0] foo0;
  output [1:0] foo1;
endmodule
