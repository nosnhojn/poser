module module2(bar, star, far, do, who, foo);
  input [1:0] bar;
  input [`BAG-1:1] star;
  input far;
  output [9:1] do;
  output [GUY:3] who;
  output foo;
endmodule
