module module3 (
  input [1:0] bar,
  input [`BAG-1:1] star,

  output [ 9 : 1]do,
  output[GUY:3]who,

  output foo,
  input far);
endmodule
