module module1(bar, foo);
  input bar;
  output foo;
endmodule
