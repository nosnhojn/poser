module module1 (
  input bar,
  output wire foo
);
endmodule
