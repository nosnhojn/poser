module module0(bar, foo);
  input bar;
  output reg foo;
endmodule
